library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all; -- Para funciones matemáticas como cos


entity Cos_LUT is
	generic(g_LUT:integer:=8
				;g_bits:integer:=32);
	port(i_angle	:	in		std_logic_vector(g_LUT-1 downto 0)
			;o_Cos	:	out	std_logic_vector(g_bits-1 downto 0)
			);
end Cos_LUT;

Architecture rtl of Cos_LUT is

	constant PI : real :=3.14159265358979323846;
	
	type t_LUT is array (0 to 2**g_LUT-1) of std_logic_vector(g_bits-1 downto 0);
	
	constant cosine_lut : t_LUT := (std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(0)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(1)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(2)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(3)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(4)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(5)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(6)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(7)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(8)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(9)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(10)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(11)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(12)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(13)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(14)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(15)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(16)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(17)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(18)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(19)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(20)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(21)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(22)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(23)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(24)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(25)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(26)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(27)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(28)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(29)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(30)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(31)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(32)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(33)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(34)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(35)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(36)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(37)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(38)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(39)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(40)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(41)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(42)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(43)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(44)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(45)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(46)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(47)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(48)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(49)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(50)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(51)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(52)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(53)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(54)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(55)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(56)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(57)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(58)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(59)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(60)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(61)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(62)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(63)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(64)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(65)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(66)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(67)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(68)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(69)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(70)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(71)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(72)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(73)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(74)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(75)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(76)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(77)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(78)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(79)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(80)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(81)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(82)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(83)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(84)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(85)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(86)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(87)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(88)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(89)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(90)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(91)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(92)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(93)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(94)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(95)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(96)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(97)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(98)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(99)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(100)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(101)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(102)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(103)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(104)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(105)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(106)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(107)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(108)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(109)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(110)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(111)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(112)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(113)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(114)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(115)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(116)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(117)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(118)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(119)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(120)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(121)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(122)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(123)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(124)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(125)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(126)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(127)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(128)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(129)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(130)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(131)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(132)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(133)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(134)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(135)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(136)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(137)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(138)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(139)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(140)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(141)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(142)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(143)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(144)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(145)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(146)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(147)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(148)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(149)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(150)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(151)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(152)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(153)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(154)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(155)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(156)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(157)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(158)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(159)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(160)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(161)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(162)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(163)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(164)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(165)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(166)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(167)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(168)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(169)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(170)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(171)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(172)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(173)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(174)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(175)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(176)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(177)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(178)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(179)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(180)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(181)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(182)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(183)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(184)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(185)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(186)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(187)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(188)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(189)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(190)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(191)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(192)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(193)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(194)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(195)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(196)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(197)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(198)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(199)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(200)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(201)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(202)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(203)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(204)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(205)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(206)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(207)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(208)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(209)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(210)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(211)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(212)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(213)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(214)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(215)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(216)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(217)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(218)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(219)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(220)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(221)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(222)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(223)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(224)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(225)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(226)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(227)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(228)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(229)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(230)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(231)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(232)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(233)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(234)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(235)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(236)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(237)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(238)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(239)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(240)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(241)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(242)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(243)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(244)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(245)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(246)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(247)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(248)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(249)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(250)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(251)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(252)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(253)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(254)/real(2**g_LUT))*PI))),g_bits)),
												std_logic_vector(to_signed(integer(floor(real(2**(g_bits-1)-1)*cos((real(255)/real(2**g_LUT))*PI))),g_bits))
	
	);

begin
	o_Cos <= cosine_LUT(to_integer(unsigned(i_angle)));
end rtl;